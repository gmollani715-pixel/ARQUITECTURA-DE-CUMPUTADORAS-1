module OR_gate{

    input wire A, //entrada A
    input wire B, //entrada B
    output wire Y //salida Y
);
    assign Y = A | B; //Operación OR
endmodule   